// module decleration.
module fun(input a,b,output y);
 //(Identifiers in this module are
 //fun (name given to the module), inputs a,b, output y and gatenames A and O
// all indentfier provided from the user side.) 
  
  and A (y,a,b);  // gate level design 
  or O (y,a,b);
  
endmodule // endmodule.

